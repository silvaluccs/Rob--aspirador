module segEeG(outSegE, outSegG);
  output outSegE, outSegG;
  
  assign outSegG = 1'b0;
  assign outSegE = 1'b0;

endmodule